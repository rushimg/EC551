`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:29:54 10/12/2012 
// Design Name: 
// Module Name:    Lab2_top 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Lab2_top(
	output [6:0] sevseg_disp,
	output [3:0] sevseg_anode,
	input	[2:0] a, b, func,
	input clk, rst, 
    );


endmodule
